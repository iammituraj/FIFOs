/*=================================================================================================================================================================================
   Design       : Dual-port RAM

   Description  : Fully synthesisable and configurable Dual-port RAM. One write port & read port.
                  - Infers Dual port Distributed RAM on FPGA Synthesisers.
                  - Configurable Data width.
                  - Configurable Depth.
                  
   Developer    : Mitu Raj, iammituraj@gmail.com
   Date         : Feb-17-2021
=================================================================================================================================================================================*/
/*=================================================================================================================================================================================
                                                                        D U A L   P O R T   R A M
=================================================================================================================================================================================*/

module my_ram   #(
                    /* Global Parameters */
                    parameter DATA_W           = 8                    ,        // Data width
                    parameter DEPTH            = 8                    ,        // Depth

                    /* Dependent Parameters */
                    parameter ADDR_W           = $clog2 (DEPTH)                // Address width 
                 )

                 (
                    /* Global */                  
                    input  logic                  clk                 ,        // Clock

                    /* Control */
                    input  logic                  i_ramen             ,        // RAM enable 
                                       
                    /* Write Port*/
                    input  logic                  i_wren              ,        // Write Enable
                    input  logic [ADDR_W - 1 : 0] i_waddr             ,        // Write-address                    
                    input  logic [DATA_W - 1 : 0] i_wdata             ,        // Write-data 
                    
                    /* Read Port */
                    input  logic [ADDR_W - 1 : 0] i_raddr             ,        // Read-address                   
                    output logic [DATA_W - 1 : 0] o_rdata                      // Read-data                   
                 );


/*---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
   Internal Registers/Signals
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*/
(* ram_style ="distributed" *)
logic [DATA_W - 1 : 0] data_rg [DEPTH] ;        // Data array


/*---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
   Synchronous logic to write to RAM
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*/
always @ (posedge clk) begin
              
   if (i_ramen) begin

      if (i_wren) begin                          
         
         data_rg [i_waddr] <= i_wdata  ;      

      end

   end

end


/*---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
   Asynchronous logic to read from RAM
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*/
assign o_rdata = data_rg [i_raddr] ;


endmodule

/*=================================================================================================================================================================================
                                                                        D U A L   P O R T   R A M
=================================================================================================================================================================================*/
